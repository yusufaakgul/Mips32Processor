library verilog;
use verilog.vl_types.all;
entity comparator32_testbench is
end comparator32_testbench;
