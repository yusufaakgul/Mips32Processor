library verilog;
use verilog.vl_types.all;
entity sign_extender_testbench is
end sign_extender_testbench;
