library verilog;
use verilog.vl_types.all;
entity shift_left2_testbench is
end shift_left2_testbench;
