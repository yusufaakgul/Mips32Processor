library verilog;
use verilog.vl_types.all;
entity alu32_testbench is
end alu32_testbench;
