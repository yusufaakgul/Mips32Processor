library verilog;
use verilog.vl_types.all;
entity mips32 is
    port(
        clk             : in     vl_logic
    );
end mips32;
