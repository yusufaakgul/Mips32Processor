library verilog;
use verilog.vl_types.all;
entity instruction_memory is
    port(
        ins             : out    vl_logic_vector(31 downto 0);
        address         : in     vl_logic_vector(11 downto 0)
    );
end instruction_memory;
