library verilog;
use verilog.vl_types.all;
entity comparator32_sign_testbench is
end comparator32_sign_testbench;
