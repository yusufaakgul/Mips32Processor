module mux32 (A,B,S,O);

input [31:0] A,B;
input S;
output [31:0] O;

mux1 mux_1 (A[0],B[0],S,O[0]),
	  mux_2 (A[1],B[1],S,O[1]),
	  mux_3 (A[2],B[2],S,O[2]),
	  mux_4 (A[3],B[3],S,O[3]),
	  mux_5 (A[4],B[4],S,O[4]),
	  mux_6 (A[5],B[5],S,O[5]),
	  mux_7 (A[6],B[6],S,O[6]),
	  mux_8 (A[7],B[7],S,O[7]),
	  mux_9 (A[8],B[8],S,O[8]),
	  mux_10 (A[9],B[9],S,O[9]),
	  mux_11 (A[10],B[10],S,O[10]),
	  mux_12 (A[11],B[11],S,O[11]),
	  mux_13 (A[12],B[12],S,O[12]),
	  mux_14 (A[13],B[13],S,O[13]),
	  mux_15 (A[14],B[14],S,O[14]),
	  mux_16 (A[15],B[15],S,O[15]),
	  mux_17 (A[16],B[16],S,O[16]),
	  mux_18 (A[17],B[17],S,O[17]),
	  mux_19 (A[18],B[18],S,O[18]),
	  mux_20 (A[19],B[19],S,O[19]),
	  mux_21 (A[20],B[20],S,O[20]),
	  mux_22 (A[21],B[21],S,O[21]),
	  mux_23 (A[22],B[22],S,O[22]),
	  mux_24 (A[23],B[23],S,O[23]),
	  mux_25 (A[24],B[24],S,O[24]),
	  mux_26 (A[25],B[25],S,O[25]),
	  mux_27 (A[26],B[26],S,O[26]),
	  mux_28 (A[27],B[27],S,O[27]),
	  mux_29 (A[28],B[28],S,O[28]),
	  mux_30 (A[29],B[29],S,O[29]),
	  mux_31 (A[30],B[30],S,O[30]),
	  mux_32 (A[31],B[31],S,O[31]);
	  
endmodule