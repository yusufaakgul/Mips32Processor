library verilog;
use verilog.vl_types.all;
entity main_control_testbench is
end main_control_testbench;
