library verilog;
use verilog.vl_types.all;
entity mux32_testbench is
end mux32_testbench;
