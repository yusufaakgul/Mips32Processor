library verilog;
use verilog.vl_types.all;
entity alu_control_testbench is
end alu_control_testbench;
