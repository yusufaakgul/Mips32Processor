library verilog;
use verilog.vl_types.all;
entity add1_testbench is
end add1_testbench;
