library verilog;
use verilog.vl_types.all;
entity address_jump_testbench is
end address_jump_testbench;
