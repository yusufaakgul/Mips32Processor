library verilog;
use verilog.vl_types.all;
entity adder32_testbench is
end adder32_testbench;
