library verilog;
use verilog.vl_types.all;
entity comparator_out_select_testbench is
end comparator_out_select_testbench;
