library verilog;
use verilog.vl_types.all;
entity zeroright16_testbench is
end zeroright16_testbench;
