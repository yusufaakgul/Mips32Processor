library verilog;
use verilog.vl_types.all;
entity mux1_testbench is
end mux1_testbench;
