module sign_extender(A,O);

input[15:0] A;
output [31:0] O;

and and_1 (O[31],A[15],A[15]),
	 and_2 (O[30],A[15],A[15]),
	 and_3 (O[29],A[15],A[15]),
	 and_4 (O[28],A[15],A[15]),
	 and_5 (O[27],A[15],A[15]),
	 and_6 (O[26],A[15],A[15]),
	 and_7 (O[25],A[15],A[15]),
	 and_8 (O[24],A[15],A[15]),
	 and_9 (O[23],A[15],A[15]),
	 and_10 (O[22],A[15],A[15]),
	 and_11 (O[21],A[15],A[15]),
	 and_12 (O[20],A[15],A[15]),
	 and_13 (O[19],A[15],A[15]),
	 and_14 (O[18],A[15],A[15]),
	 and_15 (O[17],A[15],A[15]),
	 and_16 (O[16],A[15],A[15]),
	 and_17 (O[15],A[15],A[15]),
	 and_18 (O[14],A[14],A[14]),
	 and_19 (O[13],A[13],A[13]),
	 and_20 (O[12],A[12],A[12]),
	 and_21 (O[11],A[11],A[11]),
	 and_22 (O[10],A[10],A[10]),
	 and_23 (O[9],A[9],A[9]),
	 and_24 (O[8],A[8],A[8]),
	 and_25 (O[7],A[7],A[7]),
	 and_26 (O[6],A[6],A[6]),
	 and_27 (O[5],A[5],A[5]),
	 and_28 (O[4],A[4],A[4]),
	 and_29 (O[3],A[3],A[3]),
	 and_30 (O[2],A[2],A[2]),
	 and_31 (O[1],A[1],A[1]),
	 and_32 (O[0],A[0],A[0]);
					 
endmodule
