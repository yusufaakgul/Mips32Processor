library verilog;
use verilog.vl_types.all;
entity alu1_testbench is
end alu1_testbench;
